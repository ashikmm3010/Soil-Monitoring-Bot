module ColourSensorModule();

endmodule
